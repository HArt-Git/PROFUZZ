module target(clk, rst, s_axis_tdata_7, s_axis_tdata_4, prescale_15,
     prescale_14, prescale_13, prescale_11, prescale_10, prescale_9,
     prescale_8, prescale_7, prescale_6, prescale_5, prescale_4,
     prescale_3, prescale_2, prescale_0, uart_rx_inst_g5370__7410_Y,
     uart_rx_inst_g5351__1617_Y, uart_rx_inst_prescale_reg_reg_0__Q ,
     uart_rx_inst_g5221__8246_Y, uart_rx_inst_g5306__2883_Y,
     uart_rx_inst_g5215__2802_YC, uart_rx_inst_m_axis_tvalid_reg_reg_Q,
     uart_rx_inst_bit_cnt_reg_0__Q , uart_tx_inst_g5280_Y,
     uart_rx_inst_g5319__6783_Y, uart_rx_inst_g5199__5107_YC,
     uart_rx_inst_g5377__6260_Y, uart_rx_inst_g5307__2346_Y,
     uart_rx_inst_drc_bufs5450_Y, uart_tx_inst_g5340__7482_Y,
     uart_tx_inst_g5337__6131_Y, uart_tx_inst_g5377__9945_Y,
     uart_tx_inst_prescale_reg_reg_12__Q ,
     uart_tx_inst_drc_bufs5452_Y, uart_tx_inst_prescale_reg_reg_13__Q
     , uart_rx_inst_g5241__2883_Y, uart_rx_inst_g5276__2802_Y,
     uart_rx_inst_g4043__1617_Y, uart_rx_inst_g5201__6260_Y,
     uart_rx_inst_g4051__6131_Y, uart_tx_inst_g5238__9315_YS,
     uart_tx_inst_g5376_Y, uart_tx_inst_g5273__6783_YS,
     uart_rx_inst_data_reg_reg_0__Q , uart_rx_inst_drc_bufs4064_Y,
     uart_rx_inst_g4058__9945_Y, uart_rx_inst_bit_cnt_reg_3__Q ,
     uart_rx_inst_g5394_Y, uart_rx_inst_drc_bufs5444_Y,
     uart_tx_inst_g5262_Y, uart_tx_inst_g5325__4319_Y,
     uart_tx_inst_drc_bufs5444_Y, uart_tx_inst_g5408_Y,
     uart_rx_inst_g5310__7410_Y, uart_tx_inst_drc_bufs5468_Y,
     uart_rx_inst_g5382__6783_Y, uart_tx_inst_g5313__6161_Y,
     uart_tx_inst_g5271__5526_Y,
     uart_rx_inst_m_axis_tdata_reg_reg_5__Q ,
     uart_tx_inst_drc_bufs5453_Y, uart_tx_inst_g5403__5115_Y,
     uart_rx_inst_drc_bufs5415_Y, uart_rx_inst_g5293__7482_Y,
     uart_rx_inst_g5231__7482_YC, uart_tx_inst_bit_cnt_reg_0__Q ,
     uart_rx_inst_g5352__2802_Y, uart_rx_inst_g5340__7410_Y,
     uart_rx_inst_data_reg_reg_4__Q , uart_rx_inst_g5364__6161_Y,
     uart_rx_inst_g5363__4733_Y, uart_rx_inst_g4041__6783_Y,
     uart_rx_inst_busy_reg_reg_Q, uart_rx_inst_g5373_Y,
     uart_tx_inst_g5283__1705_YS, uart_rx_inst_g4044__2802_Y,
     uart_rx_inst_g5291__1881_Y, uart_tx_inst_g5221__7098_Y,
     uart_tx_inst_drc_bufs5457_Y, uart_tx_inst_g5386__6260_YC,
     uart_tx_inst_g5273__6783_YC, uart_tx_inst_g5397__8246_Y,
     uart_rx_inst_g5329__6131_Y, uart_tx_inst_g5330__1617_Y,
     uart_rx_inst_g5323__1705_Y, uart_rx_inst_drc_bufs5447_Y,
     uart_tx_inst_g5359__5526_Y, uart_tx_inst_g5341_Y,
     uart_tx_inst_g5367__7098_Y, uart_tx_inst_g5399__6131_Y,
     uart_tx_inst_g5286__5122_Y, uart_rx_inst_drc_bufs5439_Y,
     uart_tx_inst_drc_bufs5426_Y, uart_tx_inst_g5233__4733_YC,
     uart_rx_inst_drc_bufs5419_Y, uart_tx_inst_g5386__6260_YS,
     uart_tx_inst_g5352__2398_Y, uart_tx_inst_g5353__5107_Y,
     uart_tx_inst_g5250_Y, uart_tx_inst_g5332__1705_Y,
     uart_rx_inst_data_reg_reg_6__Q ,
     uart_rx_inst_m_axis_tdata_reg_reg_6__Q ,
     uart_rx_inst_g5355__8246_Y, uart_tx_inst_g5230_Y,
     uart_rx_inst_drc_bufs5435_Y, uart_tx_inst_g5333__5122_Y,
     uart_tx_inst_g5370__1881_Y, uart_tx_inst_g5324__6260_Y,
     uart_rx_inst_prescale_reg_reg_11__Q ,
     uart_rx_inst_data_reg_reg_7__Q , uart_tx_inst_g5355_Y,
     uart_rx_inst_rxd_reg_reg_Q, uart_rx_inst_g5189__1666_Y,
     uart_tx_inst_g5322__2398_Y, uart_tx_inst_prescale_reg_reg_8__Q ,
     uart_tx_inst_g5404__7482_Y, uart_tx_inst_drc_bufs5450_Y,
     uart_rx_inst_drc_bufs5425_Y, uart_rx_inst_g5391_Y,
     uart_rx_inst_prescale_reg_reg_7__Q ,
     uart_tx_inst_prescale_reg_reg_9__Q , uart_tx_inst_g5310__5115_Y,
     uart_tx_inst_g5339__5115_Y, uart_rx_inst_drc_bufs5423_Y,
     uart_rx_inst_g5400_Y, uart_rx_inst_g5217__1705_Y,
     uart_rx_inst_drc_bufs5445_Y, uart_tx_inst_g5380__1666_Y,
     uart_rx_inst_g5203__4319_YS, uart_rx_inst_g5304__9315_Y,
     uart_tx_inst_g5251__7410_Y, uart_rx_inst_g5333__4733_Y,
     uart_rx_inst_g5287__5122_Y, uart_rx_inst_g5337__2883_Y,
     uart_tx_inst_g5245_Y, uart_tx_inst_g5257_Y,
     uart_rx_inst_g5247__7410_YC, uart_tx_inst_g5253__6417_YC,
     uart_tx_inst_g5246__2346_Y, uart_rx_inst_g5390_Y,
     uart_rx_inst_g5252__6417_Y, uart_rx_inst_g5209__6783_Y,
     uart_tx_inst_g5315__9945_Y, uart_rx_inst_prescale_reg_reg_6__Q ,
     uart_tx_inst_g5363__2802_Y, uart_rx_inst_g5378__4319_Y,
     uart_rx_inst_g5225__6131_Y, uart_tx_inst_g5242_Y,
     uart_rx_inst_prescale_reg_reg_15__Q ,
     uart_rx_inst_data_reg_reg_1__Q , uart_rx_inst_g5235__6161_YS,
     uart_tx_inst_g5358__8428_Y, uart_rx_inst_g5205__8428_Y,
     uart_tx_inst_prescale_reg_reg_16__Q , uart_rx_inst_g3770_Y,
     uart_rx_inst_drc_bufs5454_Y, uart_rx_inst_bit_cnt_reg_1__Q ,
     uart_rx_inst_g5401_Y, uart_tx_inst_g5417_Y,
     uart_tx_inst_drc_bufs5437_Y, uart_tx_inst_g5277_Y,
     uart_tx_inst_g5236__6161_Y, uart_tx_inst_g5231__7482_Y,
     uart_tx_inst_g5369_Y, uart_tx_inst_drc_bufs5440_Y,
     uart_tx_inst_prescale_reg_reg_0__Q , uart_tx_inst_g5416_Y,
     uart_rx_inst_g4053__5115_Y, uart_rx_inst_g4056__6161_Y,
     uart_rx_inst_g4049__8246_Y, uart_tx_inst_prescale_reg_reg_5__Q ,
     uart_rx_inst_g5346__4319_Y, uart_rx_inst_drc_bufs5433_Y,
     uart_tx_inst_g5215__1705_Y, uart_tx_inst_g5211_Y,
     uart_tx_inst_g5383__5477_Y, uart_tx_inst_prescale_reg_reg_15__Q ,
     uart_rx_inst_g5387_Y, uart_rx_inst_drc_bufs5453_Y,
     uart_tx_inst_g5316__2883_Y, uart_tx_inst_g5390__6783_Y,
     uart_tx_inst_g5410_Y, uart_tx_inst_drc_bufs5443_Y,
     uart_tx_inst_g5223__6131_YC, uart_rx_inst_g5246_Y,
     uart_rx_inst_g5324__5122_Y, uart_tx_inst_g5328__6783_Y,
     uart_rx_inst_prescale_reg_reg_5__Q , uart_tx_inst_g5385__5107_Y,
     s_axis_tready, m_axis_tdata_7, m_axis_tdata_3, m_axis_tdata_2,
     m_axis_tdata_1, m_axis_tdata_0, txd, rx_frame_error,
     uart_rx_inst_drc_bufs5437_A, uart_rx_inst_g5363__4733_B,
     uart_rx_inst_g5387_A, uart_rx_inst_g4044__2802_A,
     uart_rx_inst_g5210_A, uart_tx_inst_g5358__8428_C,
     uart_rx_inst_g5191__7410_B, uart_rx_inst_g5194_A,
     uart_rx_inst_g5363__4733_A, uart_rx_inst_drc_bufs5423_A,
     uart_rx_inst_data_reg_reg_3__D , uart_rx_inst_g5203__4319_B,
     uart_rx_inst_data_reg_reg_4__D , uart_tx_inst_drc_bufs5461_A,
     uart_rx_inst_g5394_A, uart_rx_inst_g5401_A,
     uart_rx_inst_drc_bufs4064_A, uart_rx_inst_g5390_A,
     uart_tx_inst_g5236__6161_A, uart_tx_inst_g5369_A,
     uart_tx_inst_g5271__5526_A, uart_rx_inst_g5334__6161_B,
     uart_rx_inst_g5364__6161_B, uart_tx_inst_g5318__1666_B,
     uart_tx_inst_data_reg_reg_6__D ,
     uart_rx_inst_m_axis_tvalid_reg_reg_D,
     uart_tx_inst_prescale_reg_reg_7__D , uart_rx_inst_g5259__8428_A,
     uart_tx_inst_g5331__2802_C, uart_tx_inst_g5263__6260_A,
     uart_rx_inst_g5332__7482_B, uart_tx_inst_g5339__5115_D,
     uart_rx_inst_g5247__7410_B, uart_rx_inst_g5226_A,
     uart_rx_inst_drc_bufs5415_A, uart_tx_inst_g5360__6783_B,
     uart_rx_inst_g5315__6260_A, uart_rx_inst_drc_bufs5450_A,
     uart_rx_inst_g5252__6417_A, uart_rx_inst_g5205__8428_A,
     uart_rx_inst_drc_bufs5434_A, uart_tx_inst_g5281__2802_A,
     uart_rx_inst_bit_cnt_reg_1__D ,
     uart_rx_inst_overrun_error_reg_reg_D,
     uart_tx_inst_prescale_reg_reg_9__D ,
     uart_rx_inst_data_reg_reg_7__D , uart_tx_inst_g5283__1705_B,
     uart_tx_inst_g5263__6260_B, uart_tx_inst_g5267_A,
     uart_tx_inst_g5316__2883_C, uart_rx_inst_bit_cnt_reg_0__D ,
     uart_tx_inst_g5278__1617_A, uart_tx_inst_drc_bufs5444_A,
     uart_rx_inst_g5305__9945_A, uart_tx_inst_drc_bufs5470_A,
     uart_tx_inst_g5223__6131_B, uart_tx_inst_g5227_A,
     uart_rx_inst_g5323__1705_A, uart_tx_inst_g5316__2883_A,
     uart_rx_inst_g5247__7410_A, uart_tx_inst_prescale_reg_reg_2__D ,
     uart_tx_inst_g5401__1881_A, uart_tx_inst_g5411_A,
     uart_rx_inst_g5333__4733_B, uart_tx_inst_g5322__2398_A,
     uart_rx_inst_data_reg_reg_6__D , uart_rx_inst_drc_bufs5418_A,
     uart_rx_inst_busy_reg_reg_D, uart_tx_inst_drc_bufs5437_A,
     uart_tx_inst_g5383__5477_B, uart_tx_inst_g5393__2802_A,
     uart_tx_inst_g5322__2398_B, uart_tx_inst_g5311__7482_C,
     uart_rx_inst_g5305__9945_B, uart_tx_inst_g5273__6783_A,
     uart_tx_inst_drc_bufs5445_A, uart_tx_inst_drc_bufs5453_A,
     uart_rx_inst_g5377__6260_A, uart_rx_inst_g5287__5122_B,
     uart_rx_inst_g5290__6131_B, uart_tx_inst_g5403__5115_B,
     uart_tx_inst_drc_bufs5440_A, uart_tx_inst_g5325__4319_B,
     uart_tx_inst_drc_bufs5434_A, uart_tx_inst_g5405_A,
     uart_tx_inst_g5367__7098_B, uart_tx_inst_g5380__1666_A,
     uart_tx_inst_g5315__9945_B, uart_rx_inst_g5231__7482_A,
     uart_rx_inst_drc_bufs5435_A, uart_rx_inst_g4049__8246_A,
     uart_tx_inst_g5286__5122_B, uart_rx_inst_g4043__1617_B,
     uart_rx_inst_g5201__6260_A, uart_tx_inst_prescale_reg_reg_8__D ,
     uart_rx_inst_g5215__2802_B, uart_rx_inst_g5218_A,
     uart_tx_inst_g5250_A, uart_rx_inst_m_axis_tdata_reg_reg_6__D ,
     uart_tx_inst_g5333__5122_A, uart_tx_inst_g5233__4733_A,
     uart_tx_inst_drc_bufs5457_A, uart_tx_inst_drc_bufs5422_A,
     uart_rx_inst_g5239__9945_B, uart_tx_inst_g5247_A,
     uart_tx_inst_g5215__1705_A, uart_tx_inst_g5245_A,
     uart_rx_inst_g5203__4319_A, uart_tx_inst_g5238__9315_A,
     uart_rx_inst_g5337__2883_C, uart_rx_inst_g3770_A,
     uart_rx_inst_g4048__5122_A, uart_tx_inst_g5328__6783_C,
     uart_rx_inst_g5307__2346_B, uart_rx_inst_g5310__7410_B,
     uart_rx_inst_g5391_A, uart_rx_inst_g5241__2883_A,
     uart_tx_inst_drc_bufs5463_A, uart_rx_inst_drc_bufs5430_A,
     uart_rx_inst_g5317__8428_B, uart_tx_inst_g5238__9315_B,
     uart_tx_inst_g5242_A, uart_rx_inst_drc_bufs5448_A,
     uart_tx_inst_g5325__4319_C, uart_rx_inst_g5233__4733_A,
     uart_tx_inst_g5283__1705_A, uart_rx_inst_g4057__9315_B,
     uart_tx_inst_drc_bufs5427_A, uart_rx_inst_g5364__6161_A,
     uart_rx_inst_g5350__3680_D, uart_rx_inst_g5382__6783_A,
     uart_rx_inst_g4056__6161_A, uart_rx_inst_g5312__5477_A,
     uart_tx_inst_drc_bufs5452_A, uart_tx_inst_prescale_reg_reg_16__D
     , uart_tx_inst_drc_bufs5460_A, uart_rx_inst_g5368__2346_S,
     uart_tx_inst_g5235_A, uart_rx_inst_g5259__8428_D,
     uart_tx_inst_g5230_A, uart_rx_inst_g4041__6783_B,
     uart_tx_inst_g5355_A, uart_tx_inst_prescale_reg_reg_0__D ,
     uart_tx_inst_g5353__5107_B, uart_rx_inst_g5306__2883_B,
     uart_rx_inst_g5320__3680_A, uart_rx_inst_g5222_A,
     uart_tx_inst_g5377__9945_A, uart_rx_inst_drc_bufs5443_A,
     uart_tx_inst_g5385__5107_A, uart_rx_inst_g5320__3680_B,
     uart_rx_inst_g5304__9315_B, uart_tx_inst_g5401__1881_C,
     uart_rx_inst_g5373_A, uart_rx_inst_data_reg_reg_0__D ,
     uart_rx_inst_g5235__6161_A, uart_rx_inst_drc_bufs5416_A,
     uart_tx_inst_data_reg_reg_1__D , uart_rx_inst_g5315__6260_B,
     uart_tx_inst_g5383__5477_A);
  input clk, rst, s_axis_tdata_7, s_axis_tdata_4, prescale_15,
       prescale_14, prescale_13, prescale_11, prescale_10, prescale_9,
       prescale_8, prescale_7, prescale_6, prescale_5, prescale_4,
       prescale_3, prescale_2, prescale_0, uart_rx_inst_g5370__7410_Y,
       uart_rx_inst_g5351__1617_Y, uart_rx_inst_prescale_reg_reg_0__Q
       , uart_rx_inst_g5221__8246_Y, uart_rx_inst_g5306__2883_Y,
       uart_rx_inst_g5215__2802_YC,
       uart_rx_inst_m_axis_tvalid_reg_reg_Q,
       uart_rx_inst_bit_cnt_reg_0__Q , uart_tx_inst_g5280_Y,
       uart_rx_inst_g5319__6783_Y, uart_rx_inst_g5199__5107_YC,
       uart_rx_inst_g5377__6260_Y, uart_rx_inst_g5307__2346_Y,
       uart_rx_inst_drc_bufs5450_Y, uart_tx_inst_g5340__7482_Y,
       uart_tx_inst_g5337__6131_Y, uart_tx_inst_g5377__9945_Y,
       uart_tx_inst_prescale_reg_reg_12__Q ,
       uart_tx_inst_drc_bufs5452_Y,
       uart_tx_inst_prescale_reg_reg_13__Q ,
       uart_rx_inst_g5241__2883_Y, uart_rx_inst_g5276__2802_Y,
       uart_rx_inst_g4043__1617_Y, uart_rx_inst_g5201__6260_Y,
       uart_rx_inst_g4051__6131_Y, uart_tx_inst_g5238__9315_YS,
       uart_tx_inst_g5376_Y, uart_tx_inst_g5273__6783_YS,
       uart_rx_inst_data_reg_reg_0__Q , uart_rx_inst_drc_bufs4064_Y,
       uart_rx_inst_g4058__9945_Y, uart_rx_inst_bit_cnt_reg_3__Q ,
       uart_rx_inst_g5394_Y, uart_rx_inst_drc_bufs5444_Y,
       uart_tx_inst_g5262_Y, uart_tx_inst_g5325__4319_Y,
       uart_tx_inst_drc_bufs5444_Y, uart_tx_inst_g5408_Y,
       uart_rx_inst_g5310__7410_Y, uart_tx_inst_drc_bufs5468_Y,
       uart_rx_inst_g5382__6783_Y, uart_tx_inst_g5313__6161_Y,
       uart_tx_inst_g5271__5526_Y,
       uart_rx_inst_m_axis_tdata_reg_reg_5__Q ,
       uart_tx_inst_drc_bufs5453_Y, uart_tx_inst_g5403__5115_Y,
       uart_rx_inst_drc_bufs5415_Y, uart_rx_inst_g5293__7482_Y,
       uart_rx_inst_g5231__7482_YC, uart_tx_inst_bit_cnt_reg_0__Q ,
       uart_rx_inst_g5352__2802_Y, uart_rx_inst_g5340__7410_Y,
       uart_rx_inst_data_reg_reg_4__Q , uart_rx_inst_g5364__6161_Y,
       uart_rx_inst_g5363__4733_Y, uart_rx_inst_g4041__6783_Y,
       uart_rx_inst_busy_reg_reg_Q, uart_rx_inst_g5373_Y,
       uart_tx_inst_g5283__1705_YS, uart_rx_inst_g4044__2802_Y,
       uart_rx_inst_g5291__1881_Y, uart_tx_inst_g5221__7098_Y,
       uart_tx_inst_drc_bufs5457_Y, uart_tx_inst_g5386__6260_YC,
       uart_tx_inst_g5273__6783_YC, uart_tx_inst_g5397__8246_Y,
       uart_rx_inst_g5329__6131_Y, uart_tx_inst_g5330__1617_Y,
       uart_rx_inst_g5323__1705_Y, uart_rx_inst_drc_bufs5447_Y,
       uart_tx_inst_g5359__5526_Y, uart_tx_inst_g5341_Y,
       uart_tx_inst_g5367__7098_Y, uart_tx_inst_g5399__6131_Y,
       uart_tx_inst_g5286__5122_Y, uart_rx_inst_drc_bufs5439_Y,
       uart_tx_inst_drc_bufs5426_Y, uart_tx_inst_g5233__4733_YC,
       uart_rx_inst_drc_bufs5419_Y, uart_tx_inst_g5386__6260_YS,
       uart_tx_inst_g5352__2398_Y, uart_tx_inst_g5353__5107_Y,
       uart_tx_inst_g5250_Y, uart_tx_inst_g5332__1705_Y,
       uart_rx_inst_data_reg_reg_6__Q ,
       uart_rx_inst_m_axis_tdata_reg_reg_6__Q ,
       uart_rx_inst_g5355__8246_Y, uart_tx_inst_g5230_Y,
       uart_rx_inst_drc_bufs5435_Y, uart_tx_inst_g5333__5122_Y,
       uart_tx_inst_g5370__1881_Y, uart_tx_inst_g5324__6260_Y,
       uart_rx_inst_prescale_reg_reg_11__Q ,
       uart_rx_inst_data_reg_reg_7__Q , uart_tx_inst_g5355_Y,
       uart_rx_inst_rxd_reg_reg_Q, uart_rx_inst_g5189__1666_Y,
       uart_tx_inst_g5322__2398_Y, uart_tx_inst_prescale_reg_reg_8__Q
       , uart_tx_inst_g5404__7482_Y, uart_tx_inst_drc_bufs5450_Y,
       uart_rx_inst_drc_bufs5425_Y, uart_rx_inst_g5391_Y,
       uart_rx_inst_prescale_reg_reg_7__Q ,
       uart_tx_inst_prescale_reg_reg_9__Q ,
       uart_tx_inst_g5310__5115_Y, uart_tx_inst_g5339__5115_Y,
       uart_rx_inst_drc_bufs5423_Y, uart_rx_inst_g5400_Y,
       uart_rx_inst_g5217__1705_Y, uart_rx_inst_drc_bufs5445_Y,
       uart_tx_inst_g5380__1666_Y, uart_rx_inst_g5203__4319_YS,
       uart_rx_inst_g5304__9315_Y, uart_tx_inst_g5251__7410_Y,
       uart_rx_inst_g5333__4733_Y, uart_rx_inst_g5287__5122_Y,
       uart_rx_inst_g5337__2883_Y, uart_tx_inst_g5245_Y,
       uart_tx_inst_g5257_Y, uart_rx_inst_g5247__7410_YC,
       uart_tx_inst_g5253__6417_YC, uart_tx_inst_g5246__2346_Y,
       uart_rx_inst_g5390_Y, uart_rx_inst_g5252__6417_Y,
       uart_rx_inst_g5209__6783_Y, uart_tx_inst_g5315__9945_Y,
       uart_rx_inst_prescale_reg_reg_6__Q ,
       uart_tx_inst_g5363__2802_Y, uart_rx_inst_g5378__4319_Y,
       uart_rx_inst_g5225__6131_Y, uart_tx_inst_g5242_Y,
       uart_rx_inst_prescale_reg_reg_15__Q ,
       uart_rx_inst_data_reg_reg_1__Q , uart_rx_inst_g5235__6161_YS,
       uart_tx_inst_g5358__8428_Y, uart_rx_inst_g5205__8428_Y,
       uart_tx_inst_prescale_reg_reg_16__Q , uart_rx_inst_g3770_Y,
       uart_rx_inst_drc_bufs5454_Y, uart_rx_inst_bit_cnt_reg_1__Q ,
       uart_rx_inst_g5401_Y, uart_tx_inst_g5417_Y,
       uart_tx_inst_drc_bufs5437_Y, uart_tx_inst_g5277_Y,
       uart_tx_inst_g5236__6161_Y, uart_tx_inst_g5231__7482_Y,
       uart_tx_inst_g5369_Y, uart_tx_inst_drc_bufs5440_Y,
       uart_tx_inst_prescale_reg_reg_0__Q , uart_tx_inst_g5416_Y,
       uart_rx_inst_g4053__5115_Y, uart_rx_inst_g4056__6161_Y,
       uart_rx_inst_g4049__8246_Y, uart_tx_inst_prescale_reg_reg_5__Q
       , uart_rx_inst_g5346__4319_Y, uart_rx_inst_drc_bufs5433_Y,
       uart_tx_inst_g5215__1705_Y, uart_tx_inst_g5211_Y,
       uart_tx_inst_g5383__5477_Y, uart_tx_inst_prescale_reg_reg_15__Q
       , uart_rx_inst_g5387_Y, uart_rx_inst_drc_bufs5453_Y,
       uart_tx_inst_g5316__2883_Y, uart_tx_inst_g5390__6783_Y,
       uart_tx_inst_g5410_Y, uart_tx_inst_drc_bufs5443_Y,
       uart_tx_inst_g5223__6131_YC, uart_rx_inst_g5246_Y,
       uart_rx_inst_g5324__5122_Y, uart_tx_inst_g5328__6783_Y,
       uart_rx_inst_prescale_reg_reg_5__Q , uart_tx_inst_g5385__5107_Y;
  output s_axis_tready, m_axis_tdata_7, m_axis_tdata_3, m_axis_tdata_2,
       m_axis_tdata_1, m_axis_tdata_0, txd, rx_frame_error,
       uart_rx_inst_drc_bufs5437_A, uart_rx_inst_g5363__4733_B,
       uart_rx_inst_g5387_A, uart_rx_inst_g4044__2802_A,
       uart_rx_inst_g5210_A, uart_tx_inst_g5358__8428_C,
       uart_rx_inst_g5191__7410_B, uart_rx_inst_g5194_A,
       uart_rx_inst_g5363__4733_A, uart_rx_inst_drc_bufs5423_A,
       uart_rx_inst_data_reg_reg_3__D , uart_rx_inst_g5203__4319_B,
       uart_rx_inst_data_reg_reg_4__D , uart_tx_inst_drc_bufs5461_A,
       uart_rx_inst_g5394_A, uart_rx_inst_g5401_A,
       uart_rx_inst_drc_bufs4064_A, uart_rx_inst_g5390_A,
       uart_tx_inst_g5236__6161_A, uart_tx_inst_g5369_A,
       uart_tx_inst_g5271__5526_A, uart_rx_inst_g5334__6161_B,
       uart_rx_inst_g5364__6161_B, uart_tx_inst_g5318__1666_B,
       uart_tx_inst_data_reg_reg_6__D ,
       uart_rx_inst_m_axis_tvalid_reg_reg_D,
       uart_tx_inst_prescale_reg_reg_7__D ,
       uart_rx_inst_g5259__8428_A, uart_tx_inst_g5331__2802_C,
       uart_tx_inst_g5263__6260_A, uart_rx_inst_g5332__7482_B,
       uart_tx_inst_g5339__5115_D, uart_rx_inst_g5247__7410_B,
       uart_rx_inst_g5226_A, uart_rx_inst_drc_bufs5415_A,
       uart_tx_inst_g5360__6783_B, uart_rx_inst_g5315__6260_A,
       uart_rx_inst_drc_bufs5450_A, uart_rx_inst_g5252__6417_A,
       uart_rx_inst_g5205__8428_A, uart_rx_inst_drc_bufs5434_A,
       uart_tx_inst_g5281__2802_A, uart_rx_inst_bit_cnt_reg_1__D ,
       uart_rx_inst_overrun_error_reg_reg_D,
       uart_tx_inst_prescale_reg_reg_9__D ,
       uart_rx_inst_data_reg_reg_7__D , uart_tx_inst_g5283__1705_B,
       uart_tx_inst_g5263__6260_B, uart_tx_inst_g5267_A,
       uart_tx_inst_g5316__2883_C, uart_rx_inst_bit_cnt_reg_0__D ,
       uart_tx_inst_g5278__1617_A, uart_tx_inst_drc_bufs5444_A,
       uart_rx_inst_g5305__9945_A, uart_tx_inst_drc_bufs5470_A,
       uart_tx_inst_g5223__6131_B, uart_tx_inst_g5227_A,
       uart_rx_inst_g5323__1705_A, uart_tx_inst_g5316__2883_A,
       uart_rx_inst_g5247__7410_A, uart_tx_inst_prescale_reg_reg_2__D
       , uart_tx_inst_g5401__1881_A, uart_tx_inst_g5411_A,
       uart_rx_inst_g5333__4733_B, uart_tx_inst_g5322__2398_A,
       uart_rx_inst_data_reg_reg_6__D , uart_rx_inst_drc_bufs5418_A,
       uart_rx_inst_busy_reg_reg_D, uart_tx_inst_drc_bufs5437_A,
       uart_tx_inst_g5383__5477_B, uart_tx_inst_g5393__2802_A,
       uart_tx_inst_g5322__2398_B, uart_tx_inst_g5311__7482_C,
       uart_rx_inst_g5305__9945_B, uart_tx_inst_g5273__6783_A,
       uart_tx_inst_drc_bufs5445_A, uart_tx_inst_drc_bufs5453_A,
       uart_rx_inst_g5377__6260_A, uart_rx_inst_g5287__5122_B,
       uart_rx_inst_g5290__6131_B, uart_tx_inst_g5403__5115_B,
       uart_tx_inst_drc_bufs5440_A, uart_tx_inst_g5325__4319_B,
       uart_tx_inst_drc_bufs5434_A, uart_tx_inst_g5405_A,
       uart_tx_inst_g5367__7098_B, uart_tx_inst_g5380__1666_A,
       uart_tx_inst_g5315__9945_B, uart_rx_inst_g5231__7482_A,
       uart_rx_inst_drc_bufs5435_A, uart_rx_inst_g4049__8246_A,
       uart_tx_inst_g5286__5122_B, uart_rx_inst_g4043__1617_B,
       uart_rx_inst_g5201__6260_A, uart_tx_inst_prescale_reg_reg_8__D
       , uart_rx_inst_g5215__2802_B, uart_rx_inst_g5218_A,
       uart_tx_inst_g5250_A, uart_rx_inst_m_axis_tdata_reg_reg_6__D ,
       uart_tx_inst_g5333__5122_A, uart_tx_inst_g5233__4733_A,
       uart_tx_inst_drc_bufs5457_A, uart_tx_inst_drc_bufs5422_A,
       uart_rx_inst_g5239__9945_B, uart_tx_inst_g5247_A,
       uart_tx_inst_g5215__1705_A, uart_tx_inst_g5245_A,
       uart_rx_inst_g5203__4319_A, uart_tx_inst_g5238__9315_A,
       uart_rx_inst_g5337__2883_C, uart_rx_inst_g3770_A,
       uart_rx_inst_g4048__5122_A, uart_tx_inst_g5328__6783_C,
       uart_rx_inst_g5307__2346_B, uart_rx_inst_g5310__7410_B,
       uart_rx_inst_g5391_A, uart_rx_inst_g5241__2883_A,
       uart_tx_inst_drc_bufs5463_A, uart_rx_inst_drc_bufs5430_A,
       uart_rx_inst_g5317__8428_B, uart_tx_inst_g5238__9315_B,
       uart_tx_inst_g5242_A, uart_rx_inst_drc_bufs5448_A,
       uart_tx_inst_g5325__4319_C, uart_rx_inst_g5233__4733_A,
       uart_tx_inst_g5283__1705_A, uart_rx_inst_g4057__9315_B,
       uart_tx_inst_drc_bufs5427_A, uart_rx_inst_g5364__6161_A,
       uart_rx_inst_g5350__3680_D, uart_rx_inst_g5382__6783_A,
       uart_rx_inst_g4056__6161_A, uart_rx_inst_g5312__5477_A,
       uart_tx_inst_drc_bufs5452_A,
       uart_tx_inst_prescale_reg_reg_16__D ,
       uart_tx_inst_drc_bufs5460_A, uart_rx_inst_g5368__2346_S,
       uart_tx_inst_g5235_A, uart_rx_inst_g5259__8428_D,
       uart_tx_inst_g5230_A, uart_rx_inst_g4041__6783_B,
       uart_tx_inst_g5355_A, uart_tx_inst_prescale_reg_reg_0__D ,
       uart_tx_inst_g5353__5107_B, uart_rx_inst_g5306__2883_B,
       uart_rx_inst_g5320__3680_A, uart_rx_inst_g5222_A,
       uart_tx_inst_g5377__9945_A, uart_rx_inst_drc_bufs5443_A,
       uart_tx_inst_g5385__5107_A, uart_rx_inst_g5320__3680_B,
       uart_rx_inst_g5304__9315_B, uart_tx_inst_g5401__1881_C,
       uart_rx_inst_g5373_A, uart_rx_inst_data_reg_reg_0__D ,
       uart_rx_inst_g5235__6161_A, uart_rx_inst_drc_bufs5416_A,
       uart_tx_inst_data_reg_reg_1__D , uart_rx_inst_g5315__6260_B,
       uart_tx_inst_g5383__5477_A;
  wire uart_rx_inst_n_1, uart_rx_inst_n_2, uart_rx_inst_n_4,
       uart_rx_inst_n_7, uart_rx_inst_n_17, uart_rx_inst_n_26,
       uart_rx_inst_n_29, uart_rx_inst_n_31;
  wire uart_rx_inst_n_33, uart_rx_inst_n_39, uart_rx_inst_n_45,
       uart_rx_inst_n_46, uart_rx_inst_n_50, uart_rx_inst_n_61,
       uart_rx_inst_n_70, uart_rx_inst_n_75;
  wire uart_rx_inst_n_83, uart_rx_inst_n_92, uart_rx_inst_n_94,
       uart_rx_inst_n_97, uart_rx_inst_n_108, uart_rx_inst_n_109,
       uart_rx_inst_n_121, uart_rx_inst_n_132;
  wire uart_rx_inst_n_139, uart_rx_inst_n_145, uart_rx_inst_n_146,
       uart_rx_inst_n_157, uart_rx_inst_n_160, uart_rx_inst_n_164,
       uart_rx_inst_n_167, uart_rx_inst_n_171;
  wire uart_rx_inst_n_174, uart_rx_inst_n_180, uart_rx_inst_n_182,
       uart_rx_inst_n_197, uart_rx_inst_n_201, uart_rx_inst_n_213,
       uart_rx_inst_n_218, uart_rx_inst_n_240;
  wire uart_rx_inst_n_241, uart_rx_inst_n_244, uart_rx_inst_n_245,
       uart_rx_inst_n_249, uart_rx_inst_n_253, uart_rx_inst_n_258,
       uart_rx_inst_n_259, uart_rx_inst_n_263;
  wire uart_rx_inst_n_266, uart_rx_inst_n_272,
       uart_rx_inst_prescale_reg17, uart_tx_inst_data_reg0,
       uart_tx_inst_n_3, uart_tx_inst_n_5, uart_tx_inst_n_10,
       uart_tx_inst_n_11;
  wire uart_tx_inst_n_15, uart_tx_inst_n_21, uart_tx_inst_n_31,
       uart_tx_inst_n_33, uart_tx_inst_n_34, uart_tx_inst_n_37,
       uart_tx_inst_n_41, uart_tx_inst_n_45;
  wire uart_tx_inst_n_46, uart_tx_inst_n_52, uart_tx_inst_n_74,
       uart_tx_inst_n_76, uart_tx_inst_n_79, uart_tx_inst_n_80,
       uart_tx_inst_n_87, uart_tx_inst_n_90;
  wire uart_tx_inst_n_96, uart_tx_inst_n_102, uart_tx_inst_n_104,
       uart_tx_inst_n_105, uart_tx_inst_n_109, uart_tx_inst_n_116,
       uart_tx_inst_n_119, uart_tx_inst_n_120;
  wire uart_tx_inst_n_121, uart_tx_inst_n_123, uart_tx_inst_n_156,
       uart_tx_inst_n_163, uart_tx_inst_n_166, uart_tx_inst_n_181,
       uart_tx_inst_n_190, uart_tx_inst_n_202;
  wire uart_tx_inst_n_232, uart_tx_inst_n_233, uart_tx_inst_n_235,
       uart_tx_inst_n_237, uart_tx_inst_prescale_reg3,
       uart_tx_inst_prescale_reg6, uart_tx_inst_prescale_reg10,
       uart_tx_inst_prescale_reg11;
  NOR2X1 uart_rx_inst_g5331__5115(.A (rst), .B
       (uart_rx_inst_g5370__7410_Y), .Y (uart_rx_inst_drc_bufs5437_A));
  BUFX2 uart_rx_inst_drc_bufs5420(.A (uart_rx_inst_g5351__1617_Y), .Y
       (uart_rx_inst_n_33));
  INVX1 uart_rx_inst_g5392(.A (uart_rx_inst_prescale_reg_reg_0__Q ),
       .Y (uart_rx_inst_g5363__4733_B));
  BUFX2 uart_tx_inst_drc_bufs5464(.A (uart_tx_inst_n_190), .Y
       (uart_tx_inst_n_5));
  DFFPOSX1 uart_rx_inst_prescale_reg_reg_9_ (.CLK (clk), .D
       (uart_rx_inst_g5221__8246_Y), .Q (uart_rx_inst_g5387_A));
  BUFX2 uart_rx_inst_drc_bufs4061(.A (uart_rx_inst_n_249), .Y
       (uart_rx_inst_g4044__2802_A));
  HAX1 uart_rx_inst_g5211__3680(.A (uart_rx_inst_g5306__2883_Y), .B
       (uart_rx_inst_g5215__2802_YC), .YC (uart_rx_inst_n_213), .YS
       (uart_rx_inst_g5210_A));
  INVX1 uart_rx_inst_g4059(.A (uart_rx_inst_m_axis_tvalid_reg_reg_Q),
       .Y (uart_rx_inst_n_245));
  OR2X1 uart_rx_inst_g5385__3680(.A (uart_rx_inst_g5364__6161_B), .B
       (uart_rx_inst_bit_cnt_reg_0__Q ), .Y (uart_rx_inst_n_70));
  DFFPOSX1 uart_tx_inst_prescale_reg_reg_4_ (.CLK (clk), .D
       (uart_tx_inst_g5280_Y), .Q (uart_tx_inst_g5358__8428_C));
  HAX1 uart_rx_inst_g5195__5477(.A (uart_rx_inst_g5319__6783_Y), .B
       (uart_rx_inst_g5199__5107_YC), .YC (uart_rx_inst_g5191__7410_B),
       .YS (uart_rx_inst_g5194_A));
  BUFX2 uart_rx_inst_drc_bufs5426(.A (uart_rx_inst_g5377__6260_Y), .Y
       (uart_rx_inst_g5363__4733_A));
  AOI22X1 uart_rx_inst_g5354__5122(.A (uart_rx_inst_g5373_A), .B
       (prescale_5), .C (prescale_4), .D (uart_rx_inst_g5350__3680_D),
       .Y (uart_rx_inst_drc_bufs5423_A));
  INVX1 uart_tx_inst_g5214(.A (uart_tx_inst_n_3), .Y
       (uart_tx_inst_n_237));
  INVX1 uart_rx_inst_g5284(.A (uart_rx_inst_n_2), .Y
       (uart_rx_inst_data_reg_reg_3__D ));
  HAX1 uart_rx_inst_g5207__5526(.A (uart_rx_inst_g5307__2346_Y), .B
       (uart_rx_inst_n_213), .YC (uart_rx_inst_g5203__4319_B), .YS
       (uart_rx_inst_n_218));
  INVX1 uart_rx_inst_g5285(.A (uart_rx_inst_drc_bufs5450_Y), .Y
       (uart_rx_inst_data_reg_reg_4__D ));
  INVX1 uart_tx_inst_g5285(.A (uart_tx_inst_n_10), .Y
       (uart_tx_inst_n_166));
  AOI22X1 uart_tx_inst_g5212__2802(.A (uart_tx_inst_n_235), .B
       (uart_tx_inst_g5340__7482_Y), .C (prescale_15), .D
       (uart_tx_inst_g5337__6131_Y), .Y (uart_tx_inst_drc_bufs5461_A));
  BUFX2 uart_tx_inst_drc_bufs5438(.A (uart_tx_inst_n_76), .Y
       (uart_tx_inst_n_31));
  AOI21X1 uart_tx_inst_g5346__2883(.A (prescale_9), .B
       (uart_tx_inst_g5377__9945_Y), .C
       (uart_tx_inst_prescale_reg_reg_12__Q ), .Y
       (uart_tx_inst_n_120));
  DFFPOSX1 uart_tx_inst_txd_reg_reg(.CLK (clk), .D
       (uart_tx_inst_drc_bufs5452_Y), .Q (txd));
  MUX2X1 uart_tx_inst_g5388__8428(.A (uart_tx_inst_g5353__5107_B), .B
       (uart_tx_inst_n_74), .S (s_axis_tready), .Y (uart_tx_inst_n_80));
  AOI22X1 uart_rx_inst_g5341__6417(.A (uart_rx_inst_g5373_A), .B
       (prescale_15), .C (prescale_14), .D
       (uart_rx_inst_g5350__3680_D), .Y (uart_rx_inst_n_109));
  AOI21X1 uart_tx_inst_g5347__2346(.A (prescale_10), .B
       (uart_tx_inst_g5377__9945_Y), .C
       (uart_tx_inst_prescale_reg_reg_13__Q ), .Y
       (uart_tx_inst_n_119));
  DFFPOSX1 uart_rx_inst_prescale_reg_reg_4_ (.CLK (clk), .D
       (uart_rx_inst_g5241__2883_Y), .Q (uart_rx_inst_g5394_A));
  DFFPOSX1 uart_rx_inst_prescale_reg_reg_1_ (.CLK (clk), .D
       (uart_rx_inst_g5276__2802_Y), .Q (uart_rx_inst_g5401_A));
  NOR2X1 uart_rx_inst_g4035__2398(.A (uart_rx_inst_g4043__1617_Y), .B
       (uart_rx_inst_n_266), .Y (uart_rx_inst_drc_bufs4064_A));
  AOI21X1 uart_tx_inst_g5343__6161(.A (prescale_11), .B
       (uart_tx_inst_g5377__9945_Y), .C (uart_tx_inst_g5383__5477_B),
       .Y (uart_tx_inst_n_123));
  DFFPOSX1 uart_rx_inst_prescale_reg_reg_14_ (.CLK (clk), .D
       (uart_rx_inst_g5201__6260_Y), .Q (uart_rx_inst_g5390_A));
  BUFX2 uart_rx_inst_drc_bufs4062(.A (uart_rx_inst_g4051__6131_Y), .Y
       (uart_rx_inst_n_241));
  INVX1 uart_tx_inst_g5237(.A (uart_tx_inst_g5238__9315_YS), .Y
       (uart_tx_inst_g5236__6161_A));
  OR2X1 uart_tx_inst_g5372__7482(.A (uart_tx_inst_g5376_Y), .B (rst),
       .Y (uart_tx_inst_g5369_A));
  INVX1 uart_tx_inst_g5272(.A (uart_tx_inst_g5273__6783_YS), .Y
       (uart_tx_inst_g5271__5526_A));
  MUX2X1 uart_rx_inst_g5358__7098(.A (uart_rx_inst_data_reg_reg_0__Q
       ), .B (m_axis_tdata_0), .S (uart_rx_inst_g5368__2346_S), .Y
       (uart_rx_inst_g5334__6161_B));
  INVX1 uart_tx_inst_g5415(.A (uart_tx_inst_g5325__4319_C), .Y
       (uart_tx_inst_n_52));
  DFFPOSX1 uart_rx_inst_frame_error_reg_reg(.CLK (clk), .D
       (uart_rx_inst_drc_bufs4064_Y), .Q (rx_frame_error));
  BUFX2 uart_tx_inst_drc_bufs5428(.A (uart_tx_inst_n_116), .Y
       (uart_tx_inst_n_41));
  OR2X1 uart_rx_inst_g4046__1705(.A (uart_rx_inst_g4058__9945_Y), .B
       (uart_rx_inst_bit_cnt_reg_3__Q ), .Y
       (uart_rx_inst_g5364__6161_B));
  AND2X1 uart_rx_inst_g5314__5107(.A (uart_rx_inst_n_33), .B
       (uart_rx_inst_g5394_Y), .Y (uart_rx_inst_n_132));
  DFFPOSX1 uart_rx_inst_m_axis_tdata_reg_reg_7_ (.CLK (clk), .D
       (uart_rx_inst_drc_bufs5444_Y), .Q (m_axis_tdata_7));
  AOI22X1 uart_tx_inst_g5261__5107(.A (uart_tx_inst_g5262_Y), .B
       (uart_tx_inst_g5340__7482_Y), .C (prescale_5), .D
       (uart_tx_inst_g5337__6131_Y), .Y (uart_tx_inst_n_190));
  AOI22X1 uart_rx_inst_g5353__1705(.A (uart_rx_inst_g5373_A), .B
       (prescale_4), .C (prescale_3), .D (uart_rx_inst_g5350__3680_D),
       .Y (uart_rx_inst_n_97));
  BUFX2 uart_tx_inst_drc_bufs5442(.A (uart_tx_inst_g5325__4319_Y), .Y
       (uart_tx_inst_g5318__1666_B));
  DFFPOSX1 uart_tx_inst_prescale_reg_reg_3_ (.CLK (clk), .D
       (uart_tx_inst_n_166), .Q (uart_tx_inst_prescale_reg3));
  OAI21X1 uart_tx_inst_g5312__4733(.A (uart_tx_inst_n_52), .B
       (uart_tx_inst_g5355_A), .C (uart_tx_inst_drc_bufs5444_Y), .Y
       (uart_tx_inst_n_156));
  OAI21X1 uart_tx_inst_g5314__9315(.A (uart_tx_inst_g5408_Y), .B
       (uart_tx_inst_g5355_A), .C (uart_tx_inst_n_21), .Y
       (uart_tx_inst_data_reg_reg_6__D ));
  BUFX2 uart_rx_inst_drc_bufs5442(.A (uart_rx_inst_g5310__7410_Y), .Y
       (uart_rx_inst_m_axis_tvalid_reg_reg_D));
  BUFX2 uart_rx_inst_drc_bufs5422(.A (uart_rx_inst_n_97), .Y
       (uart_rx_inst_n_31));
  INVX1 uart_tx_inst_g5265(.A (uart_tx_inst_drc_bufs5468_Y), .Y
       (uart_tx_inst_prescale_reg_reg_7__D ));
  OAI21X1 uart_rx_inst_g5279__1705(.A (uart_rx_inst_g4043__1617_B), .B
       (uart_rx_inst_g5323__1705_A), .C (uart_rx_inst_g5382__6783_Y),
       .Y (uart_rx_inst_g5259__8428_A));
  NAND2X1 uart_rx_inst_g5254__2398(.A (uart_rx_inst_n_75), .B
       (uart_rx_inst_n_167), .Y (uart_rx_inst_n_174));
  DFFPOSX1 uart_tx_inst_data_reg_reg_5_ (.CLK (clk), .D
       (uart_tx_inst_g5313__6161_Y), .Q (uart_tx_inst_g5331__2802_C));
  BUFX2 uart_tx_inst_drc_bufs5458(.A (uart_tx_inst_g5271__5526_Y), .Y
       (uart_tx_inst_n_11));
  BUFX2 uart_tx_inst_drc_bufs5433(.A (uart_tx_inst_n_102), .Y
       (uart_tx_inst_g5263__6260_A));
  MUX2X1 uart_tx_inst_g5362__1617(.A (prescale_15), .B
       (uart_tx_inst_g5401__1881_C), .S (uart_tx_inst_g5377__9945_Y),
       .Y (uart_tx_inst_n_104));
  MUX2X1 uart_rx_inst_g5366__9945(.A (uart_rx_inst_g5287__5122_B), .B
       (uart_rx_inst_m_axis_tdata_reg_reg_5__Q ), .S
       (uart_rx_inst_g5368__2346_S), .Y (uart_rx_inst_g5332__7482_B));
  DFFPOSX1 uart_tx_inst_s_axis_tready_reg_reg(.CLK (clk), .D
       (uart_tx_inst_drc_bufs5453_Y), .Q (s_axis_tready));
  AND2X1 uart_tx_inst_g5371__5115(.A (uart_tx_inst_g5377__9945_Y), .B
       (uart_tx_inst_g5403__5115_Y), .Y (uart_tx_inst_g5339__5115_D));
  HAX1 uart_rx_inst_g5257__6260(.A (uart_rx_inst_n_39), .B
       (uart_rx_inst_drc_bufs5415_Y), .YC (uart_rx_inst_g5247__7410_B),
       .YS (uart_rx_inst_n_171));
  OR2X1 uart_rx_inst_g5379__8428(.A (uart_rx_inst_n_266), .B
       (uart_rx_inst_n_70), .Y (uart_rx_inst_n_75));
  BUFX2 uart_rx_inst_drc_bufs5449(.A (uart_rx_inst_g5293__7482_Y), .Y
       (uart_rx_inst_n_4));
  HAX1 uart_rx_inst_g5227__1881(.A (uart_rx_inst_n_146), .B
       (uart_rx_inst_g5231__7482_YC), .YC (uart_rx_inst_n_197), .YS
       (uart_rx_inst_g5226_A));
  AOI21X1 uart_rx_inst_g5322__2802(.A (uart_rx_inst_n_75), .B
       (uart_rx_inst_n_94), .C (uart_rx_inst_g5401_A), .Y
       (uart_rx_inst_drc_bufs5415_A));
  INVX1 uart_tx_inst_g5414(.A (uart_tx_inst_bit_cnt_reg_0__Q ), .Y
       (uart_tx_inst_g5360__6783_B));
  BUFX2 uart_rx_inst_drc_bufs5421(.A (uart_rx_inst_g5352__2802_Y), .Y
       (uart_rx_inst_g5315__6260_A));
  AOI22X1 uart_rx_inst_g5292__5115(.A (uart_rx_inst_g5340__7410_Y), .B
       (uart_rx_inst_data_reg_reg_4__Q ), .C
       (uart_rx_inst_g5287__5122_B), .D (uart_rx_inst_g5364__6161_Y),
       .Y (uart_rx_inst_drc_bufs5450_A));
  INVX1 uart_rx_inst_g5356(.A (uart_rx_inst_g5363__4733_Y), .Y
       (uart_rx_inst_n_94));
  INVX1 uart_rx_inst_g3771(.A (uart_rx_inst_g4041__6783_Y), .Y
       (uart_rx_inst_n_263));
  INVX1 uart_rx_inst_g5256(.A (uart_rx_inst_n_171), .Y
       (uart_rx_inst_g5252__6417_A));
  INVX1 uart_rx_inst_g5206(.A (uart_rx_inst_n_218), .Y
       (uart_rx_inst_g5205__8428_A));
  NAND2X1 uart_rx_inst_g5359__6131(.A (uart_rx_inst_busy_reg_reg_Q), .B
       (uart_rx_inst_g5373_Y), .Y (uart_rx_inst_drc_bufs5434_A));
  INVX1 uart_tx_inst_g5282(.A (uart_tx_inst_g5283__1705_YS), .Y
       (uart_tx_inst_g5281__2802_A));
  BUFX2 uart_rx_inst_drc_bufs(.A (uart_rx_inst_g4044__2802_Y), .Y
       (uart_rx_inst_n_244));
  BUFX2 uart_rx_inst_drc_bufs5451(.A (uart_rx_inst_g5291__1881_Y), .Y
       (uart_rx_inst_n_2));
  BUFX2 uart_rx_inst_drc_bufs5440(.A (uart_rx_inst_n_174), .Y
       (uart_rx_inst_bit_cnt_reg_1__D ));
  BUFX2 uart_tx_inst_drc_bufs5454(.A (uart_tx_inst_g5221__7098_Y), .Y
       (uart_tx_inst_n_15));
  NOR3X1 uart_rx_inst_g4037__6260(.A (uart_rx_inst_n_245), .B
       (uart_rx_inst_g4041__6783_Y), .C (uart_rx_inst_g3770_A), .Y
       (uart_rx_inst_overrun_error_reg_reg_D));
  INVX1 uart_tx_inst_g5255(.A (uart_tx_inst_drc_bufs5457_Y), .Y
       (uart_tx_inst_prescale_reg_reg_9__D ));
  INVX1 uart_rx_inst_g5286(.A (uart_rx_inst_n_4), .Y
       (uart_rx_inst_data_reg_reg_7__D ));
  NOR2X1 uart_rx_inst_g4054__7482(.A (uart_rx_inst_prescale_reg17), .B
       (uart_rx_inst_g5390_A), .Y (uart_rx_inst_n_249));
  HAX1 uart_tx_inst_g5300__8246(.A (uart_tx_inst_g5386__6260_YC), .B
       (uart_tx_inst_n_34), .YC (uart_tx_inst_g5283__1705_B), .YS
       (uart_tx_inst_n_163));
  HAX1 uart_tx_inst_g5268__8428(.A (uart_tx_inst_n_37), .B
       (uart_tx_inst_g5273__6783_YC), .YC (uart_tx_inst_g5263__6260_B),
       .YS (uart_tx_inst_g5267_A));
  NOR3X1 uart_tx_inst_g5375__9315(.A (uart_tx_inst_g5403__5115_B), .B
       (uart_tx_inst_bit_cnt_reg_0__Q ), .C (uart_tx_inst_g5376_Y), .Y
       (uart_tx_inst_n_96));
  INVX1 uart_tx_inst_g5394(.A (uart_tx_inst_g5397__8246_Y), .Y
       (uart_tx_inst_n_74));
  BUFX2 uart_rx_inst_drc_bufs5436(.A (uart_rx_inst_g5329__6131_Y), .Y
       (uart_rx_inst_n_17));
  BUFX2 uart_tx_inst_drc_bufs5446(.A (uart_tx_inst_g5330__1617_Y), .Y
       (uart_tx_inst_g5316__2883_C));
  OAI21X1 uart_rx_inst_g5274__3680(.A (uart_rx_inst_g4043__1617_B), .B
       (uart_rx_inst_g5382__6783_Y), .C (uart_rx_inst_g5323__1705_Y),
       .Y (uart_rx_inst_bit_cnt_reg_0__D ));
  INVX1 uart_rx_inst_g5283(.A (uart_rx_inst_drc_bufs5447_Y), .Y
       (uart_rx_inst_n_157));
  BUFX2 uart_tx_inst_drc_bufs5430(.A (uart_tx_inst_g5359__5526_Y), .Y
       (uart_tx_inst_g5278__1617_A));
  AOI22X1 uart_tx_inst_g5326__8428(.A (uart_tx_inst_g5341_Y), .B
       (s_axis_tdata_4), .C (uart_tx_inst_g5331__2802_C), .D
       (uart_tx_inst_g5367__7098_Y), .Y (uart_tx_inst_drc_bufs5444_A));
  BUFX2 uart_rx_inst_drc_bufs5429(.A (uart_rx_inst_n_108), .Y
       (uart_rx_inst_g5305__9945_A));
  NAND2X1 uart_tx_inst_g5348__1666(.A (uart_tx_inst_g5399__6131_Y), .B
       (uart_tx_inst_n_96), .Y (uart_tx_inst_drc_bufs5470_A));
  BUFX2 uart_tx_inst_drc_bufs5459(.A (uart_tx_inst_g5286__5122_Y), .Y
       (uart_tx_inst_n_10));
  DFFPOSX1 uart_rx_inst_m_axis_tdata_reg_reg_3_ (.CLK (clk), .D
       (uart_rx_inst_drc_bufs5439_Y), .Q (m_axis_tdata_3));
  HAX1 uart_tx_inst_g5228__5115(.A (uart_tx_inst_drc_bufs5426_Y), .B
       (uart_tx_inst_g5233__4733_YC), .YC (uart_tx_inst_g5223__6131_B),
       .YS (uart_tx_inst_g5227_A));
  INVX1 uart_rx_inst_g5326(.A (uart_rx_inst_g5259__8428_D), .Y
       (uart_rx_inst_g5323__1705_A));
  INVX1 uart_tx_inst_g5407(.A (uart_tx_inst_data_reg0), .Y
       (uart_tx_inst_g5316__2883_A));
  AND2X1 uart_rx_inst_g5321__1617(.A (uart_rx_inst_drc_bufs5419_Y), .B
       (uart_rx_inst_n_61), .Y (uart_rx_inst_g5247__7410_A));
  OAI21X1 uart_tx_inst_g5320__6417(.A (uart_tx_inst_g5386__6260_YS), .B
       (uart_tx_inst_g5352__2398_Y), .C (uart_tx_inst_g5353__5107_Y),
       .Y (uart_tx_inst_prescale_reg_reg_2__D ));
  DFFPOSX1 uart_tx_inst_prescale_reg_reg_17_ (.CLK (clk), .D
       (uart_tx_inst_n_237), .Q (uart_tx_inst_g5401__1881_A));
  DFFPOSX1 uart_tx_inst_prescale_reg_reg_10_ (.CLK (clk), .D
       (uart_tx_inst_g5250_Y), .Q (uart_tx_inst_prescale_reg10));
  DFFPOSX1 uart_tx_inst_data_reg_reg_8_ (.CLK (clk), .D
       (uart_tx_inst_g5332__1705_Y), .Q (uart_tx_inst_g5411_A));
  MUX2X1 uart_rx_inst_g5369__1666(.A (uart_rx_inst_data_reg_reg_6__Q
       ), .B (uart_rx_inst_m_axis_tdata_reg_reg_6__Q ), .S
       (uart_rx_inst_g5368__2346_S), .Y (uart_rx_inst_g5333__4733_B));
  BUFX2 uart_rx_inst_drc_bufs5427(.A (uart_rx_inst_n_121), .Y
       (uart_rx_inst_n_26));
  INVX1 uart_tx_inst_g5413(.A (uart_tx_inst_g5403__5115_B), .Y
       (uart_tx_inst_g5322__2398_A));
  INVX1 uart_rx_inst_g5272(.A (uart_rx_inst_n_7), .Y
       (uart_rx_inst_data_reg_reg_6__D ));
  AOI22X1 uart_rx_inst_g5348__5526(.A (uart_rx_inst_g5373_A), .B
       (prescale_8), .C (prescale_7), .D (uart_rx_inst_g5350__3680_D),
       .Y (uart_rx_inst_drc_bufs5418_A));
  AND2X1 uart_rx_inst_g5313__2398(.A (uart_rx_inst_g5355__8246_Y), .B
       (uart_rx_inst_n_45), .Y (uart_rx_inst_busy_reg_reg_D));
  NAND3X1 uart_tx_inst_g5373__4733(.A (uart_tx_inst_data_reg0), .B
       (uart_tx_inst_g5367__7098_B), .C (uart_tx_inst_g5377__9945_Y),
       .Y (uart_tx_inst_drc_bufs5437_A));
  AOI21X1 uart_tx_inst_g5361__3680(.A (prescale_3), .B
       (uart_tx_inst_g5377__9945_Y), .C (uart_tx_inst_prescale_reg6),
       .Y (uart_tx_inst_n_105));
  DFFPOSX1 uart_tx_inst_prescale_reg_reg_14_ (.CLK (clk), .D
       (uart_tx_inst_g5230_Y), .Q (uart_tx_inst_g5383__5477_B));
  DFFPOSX1 uart_rx_inst_m_axis_tdata_reg_reg_2_ (.CLK (clk), .D
       (uart_rx_inst_drc_bufs5435_Y), .Q (m_axis_tdata_2));
  DFFPOSX1 uart_tx_inst_prescale_reg_reg_6_ (.CLK (clk), .D
       (uart_tx_inst_n_181), .Q (uart_tx_inst_prescale_reg6));
  DFFPOSX1 uart_tx_inst_bit_cnt_reg_2_ (.CLK (clk), .D
       (uart_tx_inst_g5333__5122_Y), .Q (uart_tx_inst_g5393__2802_A));
  AND2X1 uart_tx_inst_g5356__6260(.A (uart_tx_inst_g5370__1881_Y), .B
       (uart_tx_inst_n_31), .Y (uart_tx_inst_g5322__2398_B));
  BUFX2 uart_tx_inst_drc_bufs5449(.A (uart_tx_inst_g5324__6260_Y), .Y
       (uart_tx_inst_g5311__7482_C));
  INVX1 uart_rx_inst_g5403(.A (uart_rx_inst_prescale_reg_reg_11__Q ),
       .Y (uart_rx_inst_g5305__9945_B));
  BUFX2 uart_tx_inst_drc_bufs5431(.A (uart_tx_inst_n_105), .Y
       (uart_tx_inst_g5273__6783_A));
  AOI22X1 uart_rx_inst_g5273__6783(.A (uart_rx_inst_g5340__7410_Y), .B
       (uart_rx_inst_data_reg_reg_6__Q ), .C
       (uart_rx_inst_data_reg_reg_7__Q ), .D
       (uart_rx_inst_g5364__6161_Y), .Y (uart_rx_inst_n_164));
  AOI22X1 uart_tx_inst_g5329__3680(.A (uart_tx_inst_g5341_Y), .B
       (s_axis_tdata_7), .C (uart_tx_inst_g5328__6783_C), .D
       (uart_tx_inst_g5355_Y), .Y (uart_tx_inst_drc_bufs5445_A));
  OR2X1 uart_rx_inst_g4036__5107(.A (uart_rx_inst_g3770_A), .B
       (uart_rx_inst_rxd_reg_reg_Q), .Y (uart_rx_inst_n_266));
  NOR2X1 uart_tx_inst_g5342__4733(.A (uart_tx_inst_n_80), .B
       (uart_tx_inst_g5369_A), .Y (uart_tx_inst_drc_bufs5453_A));
  INVX1 uart_rx_inst_g5383(.A (uart_rx_inst_n_70), .Y
       (uart_rx_inst_g5377__6260_A));
  DFFPOSX1 uart_rx_inst_data_reg_reg_5_ (.CLK (clk), .D
       (uart_rx_inst_n_160), .Q (uart_rx_inst_g5287__5122_B));
  DFFPOSX1 uart_rx_inst_prescale_reg_reg_17_ (.CLK (clk), .D
       (uart_rx_inst_g5189__1666_Y), .Q (uart_rx_inst_prescale_reg17));
  DFFPOSX1 uart_rx_inst_data_reg_reg_2_ (.CLK (clk), .D
       (uart_rx_inst_n_157), .Q (uart_rx_inst_g5290__6131_B));
  DFFPOSX1 uart_tx_inst_bit_cnt_reg_1_ (.CLK (clk), .D
       (uart_tx_inst_g5322__2398_Y), .Q (uart_tx_inst_g5403__5115_B));
  AOI21X1 uart_tx_inst_g5364__1705(.A (prescale_5), .B
       (uart_tx_inst_g5377__9945_Y), .C
       (uart_tx_inst_prescale_reg_reg_8__Q ), .Y (uart_tx_inst_n_102));
  NAND2X1 uart_tx_inst_g5398__7098(.A (uart_tx_inst_g5404__7482_Y), .B
       (uart_tx_inst_g5403__5115_Y), .Y (uart_tx_inst_drc_bufs5440_A));
  BUFX2 uart_tx_inst_drc_bufs5435(.A (uart_tx_inst_n_109), .Y
       (uart_tx_inst_n_34));
  DFFPOSX1 uart_tx_inst_data_reg_reg_3_ (.CLK (clk), .D
       (uart_tx_inst_drc_bufs5450_Y), .Q (uart_tx_inst_g5325__4319_B));
  AND2X1 uart_rx_inst_g5302__4733(.A (uart_rx_inst_drc_bufs5425_Y), .B
       (uart_rx_inst_g5391_Y), .Y (uart_rx_inst_n_146));
  NOR3X1 uart_rx_inst_g4042__3680(.A
       (uart_rx_inst_prescale_reg_reg_7__Q ), .B
       (uart_rx_inst_g5391_A), .C (uart_rx_inst_n_244), .Y
       (uart_rx_inst_n_258));
  AOI21X1 uart_tx_inst_g5365__5122(.A (prescale_6), .B
       (uart_tx_inst_g5377__9945_Y), .C
       (uart_tx_inst_prescale_reg_reg_9__Q ), .Y
       (uart_tx_inst_drc_bufs5434_A));
  DFFPOSX1 uart_tx_inst_bit_cnt_reg_3_ (.CLK (clk), .D
       (uart_tx_inst_g5310__5115_Y), .Q (uart_tx_inst_g5405_A));
  INVX1 uart_tx_inst_g5402(.A (uart_tx_inst_g5403__5115_Y), .Y
       (uart_tx_inst_g5367__7098_B));
  OR2X1 uart_tx_inst_g5381__7410(.A (uart_tx_inst_n_87), .B
       (uart_tx_inst_prescale_reg6), .Y (uart_tx_inst_g5380__1666_A));
  BUFX2 uart_tx_inst_drc_bufs5436(.A (uart_tx_inst_g5339__5115_Y), .Y
       (uart_tx_inst_n_33));
  INVX1 uart_tx_inst_g5354(.A (uart_tx_inst_g5367__7098_Y), .Y
       (uart_tx_inst_g5315__9945_B));
  AND2X1 uart_rx_inst_g5318__5526(.A (uart_rx_inst_drc_bufs5423_Y), .B
       (uart_rx_inst_g5400_Y), .Y (uart_rx_inst_g5231__7482_A));
  AOI21X1 uart_tx_inst_g5357__4319(.A (prescale_0), .B
       (uart_tx_inst_g5377__9945_Y), .C (uart_tx_inst_prescale_reg3),
       .Y (uart_tx_inst_n_109));
  NOR2X1 uart_rx_inst_g5330__1881(.A (rst), .B (uart_rx_inst_n_83), .Y
       (uart_rx_inst_drc_bufs5435_A));
  DFFPOSX1 uart_rx_inst_prescale_reg_reg_10_ (.CLK (clk), .D
       (uart_rx_inst_g5217__1705_Y), .Q (uart_rx_inst_g4049__8246_A));
  DFFPOSX1 uart_rx_inst_m_axis_tdata_reg_reg_0_ (.CLK (clk), .D
       (uart_rx_inst_drc_bufs5445_Y), .Q (m_axis_tdata_0));
  OR2X1 uart_tx_inst_g5379__2346(.A (uart_tx_inst_g5380__1666_Y), .B
       (uart_tx_inst_g5358__8428_C), .Y (uart_tx_inst_n_90));
  INVX1 uart_tx_inst_g5299(.A (uart_tx_inst_n_163), .Y
       (uart_tx_inst_g5286__5122_B));
  INVX1 uart_rx_inst_g5402(.A (uart_rx_inst_bit_cnt_reg_0__Q ), .Y
       (uart_rx_inst_g4043__1617_B));
  INVX1 uart_rx_inst_g5202(.A (uart_rx_inst_g5203__4319_YS), .Y
       (uart_rx_inst_g5201__6260_A));
  INVX1 uart_tx_inst_g5260(.A (uart_tx_inst_n_5), .Y
       (uart_tx_inst_prescale_reg_reg_8__D ));
  HAX1 uart_rx_inst_g5219__5122(.A (uart_rx_inst_g5304__9315_Y), .B
       (uart_rx_inst_n_201), .YC (uart_rx_inst_g5215__2802_B), .YS
       (uart_rx_inst_g5218_A));
  AOI21X1 uart_tx_inst_g5345__9945(.A (prescale_8), .B
       (uart_tx_inst_g5377__9945_Y), .C (uart_tx_inst_prescale_reg11),
       .Y (uart_tx_inst_n_121));
  BUFX2 uart_tx_inst_drc_bufs5455(.A (uart_tx_inst_g5251__7410_Y), .Y
       (uart_tx_inst_g5250_A));
  BUFX2 uart_rx_inst_drc_bufs5441(.A (uart_rx_inst_g5333__4733_Y), .Y
       (uart_rx_inst_m_axis_tdata_reg_reg_6__D ));
  OR2X1 uart_tx_inst_g5366__8246(.A (uart_tx_inst_n_96), .B (rst), .Y
       (uart_tx_inst_g5333__5122_A));
  BUFX2 uart_tx_inst_drc_bufs5421(.A (uart_tx_inst_n_123), .Y
       (uart_tx_inst_g5233__4733_A));
  BUFX2 uart_rx_inst_drc_bufs5452(.A (uart_rx_inst_g5287__5122_Y), .Y
       (uart_rx_inst_n_1));
  BUFX2 uart_rx_inst_drc_bufs5414(.A (uart_rx_inst_g5337__2883_Y), .Y
       (uart_rx_inst_n_39));
  DFFPOSX1 uart_tx_inst_prescale_reg_reg_11_ (.CLK (clk), .D
       (uart_tx_inst_g5245_Y), .Q (uart_tx_inst_prescale_reg11));
  AOI22X1 uart_tx_inst_g5256__5477(.A (uart_tx_inst_g5257_Y), .B
       (uart_tx_inst_g5340__7482_Y), .C (prescale_6), .D
       (uart_tx_inst_g5337__6131_Y), .Y (uart_tx_inst_drc_bufs5457_A));
  AOI21X1 uart_tx_inst_g5344__9315(.A (prescale_7), .B
       (uart_tx_inst_g5377__9945_Y), .C (uart_tx_inst_prescale_reg10),
       .Y (uart_tx_inst_drc_bufs5422_A));
  HAX1 uart_rx_inst_g5243__2346(.A (uart_rx_inst_n_132), .B
       (uart_rx_inst_g5247__7410_YC), .YC (uart_rx_inst_g5239__9945_B),
       .YS (uart_rx_inst_n_182));
  HAX1 uart_tx_inst_g5248__1666(.A (uart_tx_inst_n_46), .B
       (uart_tx_inst_g5253__6417_YC), .YC (uart_tx_inst_n_202), .YS
       (uart_tx_inst_g5247_A));
  INVX1 uart_tx_inst_g5217(.A (uart_tx_inst_n_233), .Y
       (uart_tx_inst_g5215__1705_A));
  BUFX2 uart_tx_inst_drc_bufs5469(.A (uart_tx_inst_g5246__2346_Y), .Y
       (uart_tx_inst_g5245_A));
  AND2X1 uart_rx_inst_g5308__1666(.A (uart_rx_inst_n_29), .B
       (uart_rx_inst_g5390_Y), .Y (uart_rx_inst_g5203__4319_A));
  BUFX2 uart_tx_inst_drc_bufs5425(.A (uart_tx_inst_n_119), .Y
       (uart_tx_inst_g5238__9315_A));
  DFFPOSX1 uart_rx_inst_prescale_reg_reg_2_ (.CLK (clk), .D
       (uart_rx_inst_g5252__6417_Y), .Q (uart_rx_inst_g5337__2883_C));
  OR2X1 uart_rx_inst_g4038__4319(.A (uart_rx_inst_n_272), .B (rst), .Y
       (uart_rx_inst_g3770_A));
  INVX1 uart_rx_inst_g5408(.A (uart_rx_inst_g5364__6161_B), .Y
       (uart_rx_inst_n_46));
  INVX1 uart_rx_inst_g5409(.A (rst), .Y (uart_rx_inst_n_45));
  DFFPOSX1 uart_rx_inst_prescale_reg_reg_12_ (.CLK (clk), .D
       (uart_rx_inst_g5209__6783_Y), .Q (uart_rx_inst_g4048__5122_A));
  BUFX2 uart_rx_inst_drc_bufs4063(.A (uart_rx_inst_n_259), .Y
       (uart_rx_inst_n_240));
  DFFPOSX1 uart_tx_inst_data_reg_reg_7_ (.CLK (clk), .D
       (uart_tx_inst_g5315__9945_Y), .Q (uart_tx_inst_g5328__6783_C));
  INVX1 uart_rx_inst_g5404(.A (uart_rx_inst_prescale_reg_reg_6__Q ),
       .Y (uart_rx_inst_n_50));
  BUFX2 uart_tx_inst_drc_bufs5432(.A (uart_tx_inst_g5363__2802_Y), .Y
       (uart_tx_inst_n_37));
  XNOR2X1 uart_tx_inst_g5216__5122(.A (uart_tx_inst_n_232), .B
       (uart_tx_inst_n_104), .Y (uart_tx_inst_n_235));
  INVX1 uart_rx_inst_g5309(.A (uart_rx_inst_g5323__1705_Y), .Y
       (uart_rx_inst_n_139));
  INVX1 uart_rx_inst_g5397(.A (uart_rx_inst_g4057__9315_B), .Y
       (uart_rx_inst_g5307__2346_B));
  AOI22X1 uart_rx_inst_g5327__8246(.A (uart_rx_inst_g5373_A), .B
       (prescale_7), .C (prescale_6), .D (uart_rx_inst_g5350__3680_D),
       .Y (uart_rx_inst_n_121));
  MUX2X1 uart_rx_inst_g5349__6783(.A (uart_rx_inst_g5368__2346_S), .B
       (uart_rx_inst_m_axis_tvalid_reg_reg_Q), .S
       (uart_rx_inst_g5378__4319_Y), .Y (uart_rx_inst_g5310__7410_B));
  DFFPOSX1 uart_rx_inst_prescale_reg_reg_8_ (.CLK (clk), .D
       (uart_rx_inst_g5225__6131_Y), .Q (uart_rx_inst_g5391_A));
  INVX1 uart_rx_inst_g5242(.A (uart_rx_inst_n_182), .Y
       (uart_rx_inst_g5241__2883_A));
  AOI22X1 uart_tx_inst_g5241__9945(.A (uart_tx_inst_g5242_Y), .B
       (uart_tx_inst_g5340__7482_Y), .C (prescale_9), .D
       (uart_tx_inst_g5337__6131_Y), .Y (uart_tx_inst_drc_bufs5463_A));
  BUFX2 uart_rx_inst_drc_bufs5446(.A (uart_rx_inst_n_164), .Y
       (uart_rx_inst_n_7));
  MUX2X1 uart_rx_inst_g5367__2883(.A (uart_rx_inst_g5290__6131_B), .B
       (m_axis_tdata_2), .S (uart_rx_inst_g5368__2346_S), .Y
       (uart_rx_inst_n_83));
  AOI22X1 uart_rx_inst_g5343__2398(.A (uart_rx_inst_g5373_A), .B
       (prescale_10), .C (prescale_9), .D (uart_rx_inst_g5350__3680_D),
       .Y (uart_rx_inst_drc_bufs5430_A));
  INVX1 uart_rx_inst_g5395(.A (uart_rx_inst_prescale_reg_reg_15__Q ),
       .Y (uart_rx_inst_g5317__8428_B));
  AOI21X1 uart_tx_inst_g5351__5477(.A (prescale_14), .B
       (uart_tx_inst_g5377__9945_Y), .C (uart_tx_inst_g5401__1881_A),
       .Y (uart_tx_inst_n_116));
  HAX1 uart_tx_inst_g5243__2883(.A (uart_tx_inst_n_45), .B
       (uart_tx_inst_n_202), .YC (uart_tx_inst_g5238__9315_B), .YS
       (uart_tx_inst_g5242_A));
  AOI22X1 uart_rx_inst_g5288__8246(.A (uart_rx_inst_g5340__7410_Y), .B
       (uart_rx_inst_data_reg_reg_1__Q ), .C
       (uart_rx_inst_g5290__6131_B), .D (uart_rx_inst_g5364__6161_Y),
       .Y (uart_rx_inst_drc_bufs5448_A));
  DFFPOSX1 uart_tx_inst_data_reg_reg_4_ (.CLK (clk), .D
       (uart_tx_inst_n_156), .Q (uart_tx_inst_g5325__4319_C));
  INVX1 uart_rx_inst_g5234(.A (uart_rx_inst_g5235__6161_YS), .Y
       (uart_rx_inst_g5233__4733_A));
  BUFX2 uart_tx_inst_drc_bufs5429(.A (uart_tx_inst_g5358__8428_Y), .Y
       (uart_tx_inst_g5283__1705_A));
  DFFPOSX1 uart_rx_inst_prescale_reg_reg_13_ (.CLK (clk), .D
       (uart_rx_inst_g5205__8428_Y), .Q (uart_rx_inst_g4057__9315_B));
  AOI21X1 uart_tx_inst_g5350__6417(.A (prescale_13), .B
       (uart_tx_inst_g5377__9945_Y), .C
       (uart_tx_inst_prescale_reg_reg_16__Q ), .Y
       (uart_tx_inst_drc_bufs5427_A));
  AND2X1 uart_rx_inst_g5374__5477(.A (uart_rx_inst_g3770_Y), .B
       (uart_rx_inst_drc_bufs5454_Y), .Y (uart_rx_inst_g5364__6161_A));
  AND2X1 uart_rx_inst_g5375__2398(.A (uart_rx_inst_g5382__6783_A), .B
       (uart_rx_inst_n_70), .Y (uart_rx_inst_g5350__3680_D));
  INVX1 uart_rx_inst_g5407(.A (uart_rx_inst_n_272), .Y
       (uart_rx_inst_g5382__6783_A));
  DFFPOSX1 uart_rx_inst_prescale_reg_reg_3_ (.CLK (clk), .D
       (uart_rx_inst_n_180), .Q (uart_rx_inst_g4056__6161_A));
  MUX2X1 uart_rx_inst_g5260__5526(.A (uart_rx_inst_g5259__8428_A), .B
       (uart_rx_inst_n_139), .S (uart_rx_inst_bit_cnt_reg_1__Q ), .Y
       (uart_rx_inst_n_167));
  INVX1 uart_rx_inst_g5280(.A (uart_rx_inst_n_1), .Y
       (uart_rx_inst_n_160));
  AND2X1 uart_rx_inst_g5362__7482(.A (uart_rx_inst_n_75), .B
       (uart_rx_inst_g5401_Y), .Y (uart_rx_inst_g5312__5477_A));
  NAND3X1 uart_tx_inst_g5302__6131(.A (uart_tx_inst_g5417_Y), .B
       (uart_tx_inst_drc_bufs5437_Y), .C (uart_tx_inst_n_33), .Y
       (uart_tx_inst_drc_bufs5452_A));
  INVX1 uart_tx_inst_g5220(.A (uart_tx_inst_n_15), .Y
       (uart_tx_inst_prescale_reg_reg_16__D ));
  AOI22X1 uart_tx_inst_g5276__3680(.A (uart_tx_inst_g5277_Y), .B
       (uart_tx_inst_g5340__7482_Y), .C (prescale_2), .D
       (uart_tx_inst_g5337__6131_Y), .Y (uart_tx_inst_drc_bufs5460_A));
  AND2X1 uart_rx_inst_g5386__1617(.A (uart_rx_inst_g5382__6783_A), .B
       (uart_rx_inst_n_263), .Y (uart_rx_inst_g5368__2346_S));
  BUFX2 uart_tx_inst_drc_bufs5465(.A (uart_tx_inst_g5236__6161_Y), .Y
       (uart_tx_inst_g5235_A));
  AOI22X1 uart_rx_inst_g5342__5477(.A (uart_rx_inst_g5373_A), .B
       (prescale_9), .C (prescale_8), .D (uart_rx_inst_g5350__3680_D),
       .Y (uart_rx_inst_n_108));
  OAI21X1 uart_rx_inst_g5339__1666(.A (uart_rx_inst_n_46), .B
       (uart_rx_inst_n_266), .C (uart_rx_inst_n_92), .Y
       (uart_rx_inst_g5259__8428_D));
  BUFX2 uart_tx_inst_drc_bufs5467(.A (uart_tx_inst_g5231__7482_Y), .Y
       (uart_tx_inst_g5230_A));
  INVX1 uart_tx_inst_g5270(.A (uart_tx_inst_n_11), .Y
       (uart_tx_inst_n_181));
  INVX1 uart_rx_inst_g5406(.A (uart_rx_inst_rxd_reg_reg_Q), .Y
       (uart_rx_inst_g4041__6783_B));
  INVX1 uart_rx_inst_g5357(.A (uart_rx_inst_g5364__6161_Y), .Y
       (uart_rx_inst_n_92));
  AND2X1 uart_tx_inst_g5368__6131(.A (uart_tx_inst_g5369_Y), .B
       (uart_tx_inst_drc_bufs5440_Y), .Y (uart_tx_inst_g5355_A));
  OAI21X1 uart_tx_inst_g5321__5477(.A
       (uart_tx_inst_prescale_reg_reg_0__Q ), .B
       (uart_tx_inst_g5352__2398_Y), .C (uart_tx_inst_g5353__5107_Y),
       .Y (uart_tx_inst_prescale_reg_reg_0__D ));
  OR2X1 uart_tx_inst_g5391__3680(.A (uart_tx_inst_g5397__8246_Y), .B
       (uart_tx_inst_g5416_Y), .Y (uart_tx_inst_g5353__5107_B));
  OR2X1 uart_rx_inst_g4050__7098(.A (uart_rx_inst_g4053__5115_Y), .B
       (uart_rx_inst_g4056__6161_Y), .Y (uart_rx_inst_n_253));
  INVX1 uart_rx_inst_g5389(.A (uart_rx_inst_g4048__5122_A), .Y
       (uart_rx_inst_g5306__2883_B));
  BUFX2 uart_rx_inst_drc_bufs5428(.A (uart_rx_inst_n_109), .Y
       (uart_rx_inst_g5320__3680_A));
  HAX1 uart_rx_inst_g5223__7098(.A (uart_rx_inst_n_145), .B
       (uart_rx_inst_n_197), .YC (uart_rx_inst_n_201), .YS
       (uart_rx_inst_g5222_A));
  NAND3X1 uart_rx_inst_g4040__5526(.A (uart_rx_inst_n_241), .B
       (uart_rx_inst_g4049__8246_Y), .C (uart_rx_inst_n_258), .Y
       (uart_rx_inst_n_259));
  NOR3X1 uart_tx_inst_g5378__2883(.A (uart_tx_inst_prescale_reg3), .B
       (uart_tx_inst_prescale_reg_reg_5__Q ), .C (uart_tx_inst_n_90),
       .Y (uart_tx_inst_g5377__9945_A));
  BUFX2 uart_rx_inst_drc_bufs5424(.A (uart_rx_inst_g5346__4319_Y), .Y
       (uart_rx_inst_n_29));
  NAND2X1 uart_rx_inst_g5253__5477(.A (uart_rx_inst_n_75), .B
       (uart_rx_inst_drc_bufs5433_Y), .Y (uart_rx_inst_drc_bufs5443_A));
  BUFX2 uart_tx_inst_drc_bufs5466(.A (uart_tx_inst_g5215__1705_Y), .Y
       (uart_tx_inst_n_3));
  OR2X1 uart_tx_inst_g5387__4319(.A (uart_tx_inst_n_79), .B
       (uart_tx_inst_prescale_reg10), .Y (uart_tx_inst_g5385__5107_A));
  INVX1 uart_rx_inst_g5393(.A (uart_rx_inst_g4056__6161_A), .Y
       (uart_rx_inst_n_61));
  INVX1 uart_rx_inst_g5399(.A (uart_rx_inst_prescale_reg17), .Y
       (uart_rx_inst_g5320__3680_B));
  INVX1 uart_rx_inst_g5396(.A (uart_rx_inst_g4049__8246_A), .Y
       (uart_rx_inst_g5304__9315_B));
  DFFPOSX1 uart_tx_inst_prescale_reg_reg_18_ (.CLK (clk), .D
       (uart_tx_inst_g5211_Y), .Q (uart_tx_inst_g5401__1881_C));
  DFFPOSX1 uart_rx_inst_m_axis_tdata_reg_reg_1_ (.CLK (clk), .D
       (uart_rx_inst_n_17), .Q (m_axis_tdata_1));
  OR2X1 uart_tx_inst_g5382__6417(.A (uart_tx_inst_g5383__5477_Y), .B
       (uart_tx_inst_prescale_reg_reg_15__Q ), .Y (uart_tx_inst_n_87));
  AND2X1 uart_rx_inst_g5376__5107(.A (uart_rx_inst_g5382__6783_A), .B
       (uart_rx_inst_g5377__6260_A), .Y (uart_rx_inst_g5373_A));
  BUFX2 uart_tx_inst_drc_bufs5424(.A (uart_tx_inst_n_120), .Y
       (uart_tx_inst_n_45));
  OR2X1 uart_rx_inst_g4039__8428(.A (uart_rx_inst_n_240), .B
       (uart_rx_inst_n_253), .Y (uart_rx_inst_n_272));
  AND2X1 uart_rx_inst_g5303__6161(.A (uart_rx_inst_n_26), .B
       (uart_rx_inst_g5387_Y), .Y (uart_rx_inst_n_145));
  INVX1 uart_rx_inst_g5282(.A (uart_rx_inst_drc_bufs5453_Y), .Y
       (uart_rx_inst_data_reg_reg_0__D ));
  AND2X1 uart_rx_inst_g5316__4319(.A (uart_rx_inst_n_31), .B
       (uart_rx_inst_n_50), .Y (uart_rx_inst_g5235__6161_A));
  AOI22X1 uart_rx_inst_g5365__9315(.A (uart_rx_inst_g5364__6161_B), .B
       (uart_rx_inst_drc_bufs5454_Y), .C (uart_rx_inst_g4041__6783_B),
       .D (uart_rx_inst_g4043__1617_Y), .Y
       (uart_rx_inst_drc_bufs5416_A));
  DFFPOSX1 uart_tx_inst_data_reg_reg_0_ (.CLK (clk), .D
       (uart_tx_inst_g5316__2883_Y), .Q (uart_tx_inst_data_reg0));
  OR2X1 uart_tx_inst_g5389__5526(.A (uart_tx_inst_g5390__6783_Y), .B
       (uart_tx_inst_prescale_reg11), .Y (uart_tx_inst_n_79));
  OAI21X1 uart_tx_inst_g5317__2346(.A (uart_tx_inst_g5410_Y), .B
       (uart_tx_inst_g5315__9945_B), .C (uart_tx_inst_drc_bufs5443_Y),
       .Y (uart_tx_inst_data_reg_reg_1__D ));
  HAX1 uart_tx_inst_g5218__8246(.A (uart_tx_inst_n_41), .B
       (uart_tx_inst_g5223__6131_YC), .YC (uart_tx_inst_n_232), .YS
       (uart_tx_inst_n_233));
  AND2X1 uart_rx_inst_g5245__1666(.A (uart_rx_inst_g5246_Y), .B
       (uart_rx_inst_g5324__5122_Y), .Y (uart_rx_inst_n_180));
  BUFX2 uart_tx_inst_drc_bufs5448(.A (uart_tx_inst_g5328__6783_Y), .Y
       (uart_tx_inst_n_21));
  BUFX2 uart_tx_inst_drc_bufs5423(.A (uart_tx_inst_n_121), .Y
       (uart_tx_inst_n_46));
  NAND2X1 uart_tx_inst_g5392__1617(.A (uart_tx_inst_bit_cnt_reg_0__Q
       ), .B (uart_tx_inst_g5399__6131_Y), .Y (uart_tx_inst_n_76));
  INVX1 uart_rx_inst_g5398(.A (uart_rx_inst_prescale_reg_reg_5__Q ),
       .Y (uart_rx_inst_g5315__6260_B));
  OR2X1 uart_tx_inst_g5384__2398(.A (uart_tx_inst_g5385__5107_Y), .B
       (uart_tx_inst_prescale_reg_reg_13__Q ), .Y
       (uart_tx_inst_g5383__5477_A));
endmodule
